library ieee;
use ieee.std_logic_1164.all;

entity Transmitter is
port(data: in std_logic_vector (7 downto 0);
clk,parity_type,go: in std_logic;
txd, txrdy, txe: out std_logic);
end;

architecture one of Transmitter is

component generator
generic(N:  integer:= 50000000;
		  DC: integer:= 25000000);
port(
clkin: in std_logic;
clkout: buffer std_logic:='1');
end component;

component PISO
generic (n:integer:=4);
port(data: std_logic_vector (n-1 downto 0);
clk,sel: in std_logic;
Q,txe,txrdy:out std_logic);
end component;

component parity_gen
generic (N: integer:=4);
port(
inpt: std_logic_vector(N-1 downto 0);
outpt: out std_logic);
end component;

signal Parity,outxor,internclk: std_logic;
signal sdata: std_logic_vector(10 downto 0);

begin
sdata <= '1' & Parity & data & '0';
U1: PISO generic map (11) port map (sdata, internclk, go, txd, txe, txrdy);
U2: Generator generic map (5208,2604) port map (clk, internclk);
U3: Parity_Gen Generic map (8) port map (data,outxor);
Parity <= '1' when (parity_type = '0' and outxor = '0') else '0';
end;


-- / Parity_Gen \ --
library ieee;
use ieee.std_logic_1164.all;

entity Parity_Gen is
generic (N: integer:=4);
port(
inpt: std_logic_vector(N-1 downto 0);
outpt: out std_logic);
end;

architecture one of Parity_Gen is
begin
process(inpt)
variable x: std_logic;
begin
x:='0';
for i in 0 to N-1 loop
x := x xor inpt(i);
end loop;
outpt <= x;
end process;
end;

-- / Generator \ --
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Generator is
generic(N:  integer:= 50000000;
		  DC: integer:= 25000000);
port(
clkin: in std_logic;
clkout: buffer std_logic:='1');
end;

architecture one of Generator is
signal count: integer range 0 to N := 0;
begin
process(clkin)
begin
if (clkin 'event and clkin = '1') then 
	if (count = N) then
		count <= 0;
		clkout <= '1';
	elsif (count = DC) then
		count <= count + 1;
		clkout <= '0';
	else
		count <= count + 1;
	end if;
end if;
end process;
end;

-- / PISO \ --
library ieee;
use ieee.std_logic_1164.all;

entity PISO is 
generic (n:integer:=4);
port(data: std_logic_vector (n-1 downto 0);
clk,sel: in std_logic;
Q,txe,txrdy:out std_logic);
end;

architecture one of PISO is

signal sq: std_logic_vector (n-1 downto 0);
signal stxrdy,ntxe: std_logic;
signal zvec: std_logic_vector(n-1 downto 0):= (others => '0');

begin
txrdy <= stxrdy;
process(clk)
begin
for i in 0 to n-1 loop
	if (clk='1' and clk'event) then
		if (sel='0') then
			sq <= data;
		else
			sq <= '0' & sq (n-1 downto 1);
		end if;
	end if;
end loop;

if (clk 'event and clk = '1') then
	if (data = zvec) then
		stxrdy <= '0';
	else
		stxrdy <= '1';
	end if;
end if;

end process;

q<=sq(0);
txe<= not ntxe;

process(sq)
variable x: std_logic;
begin
x:='0';
for i in 0 to n-1 loop
x:= x or sq(i);
end loop;
ntxe<=x;
end process; 

end;
