library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;

entity upcount is
port (
Clear, Clock,rst: in std_logic;
Q : out std_logic_vector(1 downto 0));
end;

architecture Behavior of upcount is

signal Count : std_logic_vector(1 downto 0);

begin
process (rst,Clock)
begin
if (rst = '0') then count <= (others => '0');
elsif (Clock 'event and Clock = '1') then
	if (Clear = '1') then
		Count <= "00";
	else
		Count <= Count + 1;
	end if;
end if;

end process;

Q <= Count;
end;

library ieee;
use ieee.std_logic_1164.all;

entity dec3to8 is
port ( W : in std_logic_vector(2 downto 0);
En : in std_logic;
Y : out std_logic_vector(0 to 7));
end;

architecture Behavior of dec3to8 is
begin

process (W, En)
begin
if (En = '1') then
	case W is
	when "000"  => Y <= "00000001";
	when "001"  => Y <= "00000010";
	when "010"  => Y <= "00000100";
	when "011"  => Y <= "00001000";
	when "100"  => Y <= "00010000";
	when "101"  => Y <= "00100000";
	when "110"  => Y <= "01000000";
	when others => Y <= "10000000";
	end case;
else
	Y <= "00000000";
end if;
end process;
end Behavior;


library ieee;
use ieee.std_logic_1164.all;

entity regn is
generic (n : integer := 16);
port (
R: in std_logic_vector(n-1 downto 0);
rst, Rin, Clock: in std_logic;
Q: buffer std_logic_vector(n-1 downto 0));
end;

architecture Behavior of regn is
begin
process (rst,Clock)
begin
if (rst = '0') then Q <= (others =>'0');
elsif (Clock 'event and Clock = '1') then
	if (Rin = '1') then
		Q <= R;
	end if;
end if;
end process;
end;


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ALU is
port(
A,B: in std_logic_vector (15 downto 0);
addsub: in std_logic;
outpt: out std_logic_vector(15 downto 0));
end;

architecture one of ALU is
begin
outpt <= A + B when addsub = '0' else A - B ;
end;


library ieee;
use ieee.std_logic_1164.all;
 
entity mux is
port( 
r0,r1,r2,r3,r4,r5,r6,r7,din,g : in std_logic_vector (15 downto 0);
gout,dout: in std_logic;
rout: in std_logic_vector (7 downto 0);
busa: out std_logic_vector (15 downto 0));
end;
 
architecture bhv of mux is
begin
process (r0,r1,r2,r3,r4,r5,r6,r7,din,g,gout,dout,rout) is
begin
	if (gout = '1') then
		busa <= g;
	elsif (dout = '1') then
		busa<=din;
	else
		case (rout) is
		when "10000000" => busa <= r7;
		when "01000000" => busa <= r6;
		when "00100000" => busa <= r5;
		when "00010000" => busa <= r4;
		when "00001000" => busa <= r3;
		when "00000100" => busa <= r2;
		when "00000010" => busa <= r1;
		when others 	 => busa <= r0;
		end case;
		end if;
end process;
end;


library ieee;
use ieee.std_logic_1164.all;

entity MPU is
port(
clk,run,reset: in std_logic;
Din: in std_logic_vector(15 downto 0);
Done: out std_logic);
end;

architecture one of MPU is

-- / Components \ --

component regn
generic (n : INTEGER := 16);
port (
R: in STD_LOGIC_VECTOR(n-1 DOWNTO 0);
rst, Rin, Clock: in STD_LOGIC;
Q: buffer STD_LOGIC_VECTOR(n-1 DOWNTO 0));
end component;

component mux
port(
r0,r1,r2,r3,r4,r5,r6,r7,din,g : in STD_LOGIC_vector (15 downto 0);
gout,dout: in STD_LOGIC;
rout: in std_logic_vector (7 downto 0);
busa: out STD_LOGIC_vector (15 downto 0));
end component;

component ALU
port(
A,B: in std_logic_vector (15 downto 0);
addsub: in std_logic;
outpt: out std_logic_vector(15 downto 0));
end component;

component upcount
port(
Clear, Clock,rst: in std_logic;
Q: out std_Logic_vector(1 DOWNTO 0));
end component;

component ControlUnit
port(
Instruction: in std_logic_vector(8 downto 0);
run,reset: in std_logic;
count: in std_logic_vector(1 downto 0);

clear,Done: buffer std_logic;
Dinout,Gout,Gin,Ain,IRin,AddSub: out std_logic;
Rin:  out std_logic_vector(7 downto 0);
Rout: out std_logic_vector(7 downto 0));
end component;

-- / Components \ --

-- / Signals \ --
signal R0,R1,R2,R3,R4,R5,R6,R7: std_logic_vector(15 downto 0);
signal Gout: std_logic_vector(15 downto 0);
signal busa: std_logic_vector(15 downto 0);
signal EnReg: std_logic_vector(7 downto 0);
signal Ain,Gin,IRin: std_logic;
signal ALUout,ALUin: std_logic_vector(15 downto 0);
signal Instruction: std_logic_vector(8 downto 0);
signal sel: std_logic_vector(7 downto 0);
signal sg,sd: std_logic;
signal selALU: std_logic;
signal count: std_logic_vector(1 downto 0);
signal clrCount: std_logic;
-- / Signals \ --

begin
-- Rx:   regn generic map (16) port map (Datain, 			 En,       clk, Q);
   Reg0: regn generic map (16) port map (busa,   			 reset, EnReg(0), clk, R0);
   Reg1: regn generic map (16) port map (busa,   			 reset, EnReg(1), clk, R1);
   Reg2: regn generic map (16) port map (busa,   			 reset, EnReg(2), clk, R2);
   Reg3: regn generic map (16) port map (busa,   			 reset, EnReg(3), clk, R3);
   Reg4: regn generic map (16) port map (busa,   			 reset, EnReg(4), clk, R4);
   Reg5: regn generic map (16) port map (busa,   			 reset, EnReg(5), clk, R5);
   Reg6: regn generic map (16) port map (busa,   			 reset, EnReg(6), clk, R6);
   Reg7: regn generic map (16) port map (busa,   			 reset, EnReg(7), clk, R7);
   G:    regn generic map (16) port map (ALUout, 			 reset, Gin,      clk, Gout);
	A:    regn generic map (16) port map (busa,            reset, Ain,      clk, ALUin);
	IR:   regn generic map (9)  port map (Din(15 downto 7), reset, IRin,     clk, Instruction);

U0: ControlUnit port map (Instruction, run, reset,count,clrCount,Done,sd,sg,Gin,Ain,IRin,selALU,EnReg,sel);
U1: upcount port map (clrCount,clk,reset,count);

MultiPlexer: mux port map (R0,R1,R2,R3,R4,R5,R6,R7,Din,Gout,sg,sd,sel,busa);
ArithLogicUnit: ALU port map (ALUin,busa,selALU,ALUout);
end;


library ieee;
use ieee.std_logic_1164.all;

entity ControlUnit is
port(

Instruction: in std_logic_vector(8 downto 0);
run,reset: in std_logic;
count: in std_logic_vector(1 downto 0);

clear,Done: buffer std_logic;
Dinout,Gout,Gin,Ain,IRin,AddSub: out std_logic;
Rin:  out std_logic_vector(7 downto 0);
Rout: out std_logic_vector(7 downto 0));

end;

architecture one of ControlUnit is

component dec3to8
port(
w:  in std_logic_vector(2 downto 0);
En: in std_logic;
y:  out std_logic_vector(0 to 7));
end component;

signal Enrun: std_logic:='0';
signal EnDecin,EnDecout: std_logic;
signal AddrRegIn:  std_logic_vector(2 downto 0);
signal AddrRegOut: std_logic_vector(2 downto 0);

begin

DecEnIn:  dec3to8 port map (AddrRegIn,  EnDecin,  Rin);
DecEnOut: dec3to8 port map (AddrRegOut, EnDecout, Rout);

clear <= Done;

process (run,Done)
begin
	if (run = '1') then Enrun <='1';
	elsif (Done = '1') then Enrun <= '0';
	else Enrun <= Enrun; end if;
end process;

--
-- |---------------------------
-- |       |\            |\   |
-- |-------|0|-----------|0|------Enrun
--   '0'---|1|     '1'---|1|
--	        |/            |/
--          |             |
--          |             |
--         Done          run



process(count,Enrun,reset)
begin

--AddrRegIn  <= Instruction(5 downto 3); -- RxIn
--AddrRegOut <= Instruction(2 downto 0); -- RyOut
--AddrRegIn  <= Instruction(2 downto 0); -- RyIn
--AddrRegOut <= Instruction(5 downto 3); -- RxOut

if (reset = '0') then Done <= '0';
elsif (Enrun = '1') then
case count is
when "00" => Done <= '0'; IRin <= '1'; -- Fetch
			 EnDecin <= '0'; EnDecout <= '0';
			 Dinout <= '0'; Gout <= '0';
			 AddSub <= '0'; Ain <= '0'; Gin <= '0';
when "01" => IRin <= '0'; -- T1
	case Instruction(8 downto 6) is
	when "000"  => EnDecin <= '1'; EnDecout <= '1';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0';
				   Done <= '1';
				   AddrRegOut <= Instruction (2 downto 0); AddrRegIn <= Instruction (5 downto 3);
	when "001"  => EnDecin <= '1'; EnDecout <= '0';
				   Dinout <= '1'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0';
				   Done <= '1'; AddrRegIn  <= Instruction(5 downto 3);
	when "010"  => EnDecin <= '0'; EnDecout <= '1';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '1'; Gin <= '0';
				   Done <= '0'; AddrRegOut <= Instruction(5 downto 3);
	when "011"  => EnDecin <= '0'; EnDecout <= '1';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '1'; Ain <= '1'; Gin <= '0';
				   Done <= '0'; AddrRegOut <= Instruction(5 downto 3);
	when others => EnDecin <= '0'; EnDecout <= '0';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0'; Done <= '0';
	end case;
when "10" => -- T2
	case Instruction(8 downto 6) is
	when "010"  => EnDecin <= '0'; EnDecout <= '1';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '1';
				   Done <= '0'; AddrRegOut <= Instruction(2 downto 0); -- Add
	when "011"  => EnDecin <= '0'; EnDecout <= '1';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '1'; Ain <= '0'; Gin <= '1';
				   Done <= '0'; AddrRegOut <= Instruction(2 downto 0); -- Sub
	when others => EnDecin <= '0'; EnDecout <= '0';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0'; Done <= '0';
	end case;
when others => Done <= '1'; -- T3
	case Instruction(8 downto 6) is
	when "010"  => EnDecin <= '1'; EnDecout <= '0';
				   Dinout <= '0'; Gout <= '1';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0';
				   AddrRegIn <= Instruction(5 downto 3); -- Add
	when "011"  => EnDecin <= '1'; EnDecout <= '0';
				   Dinout <= '0'; Gout <= '1'; 
				   AddSub <= '1'; Ain <= '0'; Gin <= '0';
				   AddrRegIn <= Instruction(5 downto 3); -- Sub
	when others => EnDecin <= '0'; EnDecout <= '0';
				   Dinout <= '0'; Gout <= '0';
				   AddSub <= '0'; Ain <= '0'; Gin <= '0';
	end case;
end case;
end if;
end process;
end;


