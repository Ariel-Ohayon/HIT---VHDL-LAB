--LIBRARY ieee; USE ieee.std_logic_1164.all;
--USE ieee.std_logic_signed.all;
--
--ENTITY proc IS
--PORT (
--DIN : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
--Resetn, Clock, Run : IN STD_LOGIC;
--Done : BUFFER STD_LOGIC;
--BusWires : BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0));
--END;
--
--ARCHITECTURE Behavior OF proc IS
--... declare components
--... declare signals
--BEGIN
--
--Clear <= ...
--Tstep: upcount PORT MAP (Clear, Clock, Tstep_Q);
--I <= IR(1 TO 3);
--decX: dec3to8 PORT MAP (IR(4 TO 6), '1', Xreg);
--decY: dec3to8 PORT MAP (IR(7 TO 9), '1', Yreg);
--
--controlsignals: PROCESS (Tstep_Q, I, Xreg, Yreg)
--BEGIN
--... specify initial values
--CASE Tstep_Q IS
--WHEN "00" => -- store DIN in IR as long as Tstep_Q = 0
--IRin <= ’1’;
--WHEN "01" => -- define signals in time step T1
--CASE I IS
--...
--END CASE;
--WHEN "10" => -- define signals in time step T2
--CASE I IS
--...
--END CASE;
--WHEN "11" => -- define signals in time step T3
--	CASE I IS
--
--	END CASE;
--END CASE;
--END PROCESS;
--reg_0: regn PORT MAP (BusWires, Rin(0), Clock, R0);
--... instantiate other registers and the adder/subtracter unit
--... define the bus
--END Behavior;